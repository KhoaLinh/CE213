library verilog;
use verilog.vl_types.all;
entity test_Squareroot is
    port(
        \out\           : out    vl_logic
    );
end test_Squareroot;
