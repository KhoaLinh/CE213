library verilog;
use verilog.vl_types.all;
entity lnx_vlg_vec_tst is
end lnx_vlg_vec_tst;
