library verilog;
use verilog.vl_types.all;
entity REG16bit_vlg_check_tst is
    port(
        reg_next        : in     vl_logic_vector(15 downto 0);
        sampler_rx      : in     vl_logic
    );
end REG16bit_vlg_check_tst;
