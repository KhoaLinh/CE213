library verilog;
use verilog.vl_types.all;
entity CAS_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        cin             : in     vl_logic;
        control         : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end CAS_vlg_sample_tst;
