library verilog;
use verilog.vl_types.all;
entity CounterCheck_vlg_vec_tst is
end CounterCheck_vlg_vec_tst;
