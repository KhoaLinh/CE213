library verilog;
use verilog.vl_types.all;
entity clock_1s_vlg_check_tst is
    port(
        clk             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end clock_1s_vlg_check_tst;
