library verilog;
use verilog.vl_types.all;
entity d_ff_struct_vlg_vec_tst is
end d_ff_struct_vlg_vec_tst;
