library verilog;
use verilog.vl_types.all;
entity MUL_vlg_vec_tst is
end MUL_vlg_vec_tst;
