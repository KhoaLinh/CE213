library verilog;
use verilog.vl_types.all;
entity Data_pipeline_Beha_vlg_vec_tst is
end Data_pipeline_Beha_vlg_vec_tst;
