module tbALU();

reg [31:0] inA;
reg [31:0] inB;
reg [2:0] s;
wire [31:0] result;
ALU alu1(result,inA,inB,s);
initial
begin
    inA = 0;
    inB = 0;
    s = 0;
    #20
    inA = 32'b00000000000000000000000000000001;
    inB = 32'b00000000000000000000000000000011;
    s = 3'b000;
    #20
    inA = 32'b00000000000000000000000000000001;
    inB = 32'b00000000000000000000000000000011;
    s = 3'b001;
    #20
    inA = 32'b00000000000000000000000000000001;
    inB = 32'b00000000000000000000000000000011;
    s = 3'b010;
    #20
    inA = 32'b00000000000000000000000000000001;
    inB = 32'b00000000000000000000000000000011;
    s = 3'b011;
    #20
    inA = 32'b00000000000000000000000000000001;
    inB = 32'b00000000000000000000000000000011;
    s = 3'b100;
    #20
    inA = 32'b00000000000000000000000000000001;
    inB = 32'b00000000000000000000000000000011;
    s = 3'b101;
    #20
    inA = 32'b00000000000000000000000000000001;
    inB = 32'b00000000000000000000000000000011;
    s = 3'b110;
    #20
    inA = 32'b00000000000000000000000000000001;
    inB = 32'b00000000000000000000000000000011;
    s = 3'b111;
    #20
    $stop;
end

endmodule