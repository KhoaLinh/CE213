library verilog;
use verilog.vl_types.all;
entity bcd_counter_vlg_vec_tst is
end bcd_counter_vlg_vec_tst;
