library verilog;
use verilog.vl_types.all;
entity clockedD_latch_vlg_vec_tst is
end clockedD_latch_vlg_vec_tst;
