library verilog;
use verilog.vl_types.all;
entity REG16bit_vlg_vec_tst is
end REG16bit_vlg_vec_tst;
