library verilog;
use verilog.vl_types.all;
entity getMode_vlg_vec_tst is
end getMode_vlg_vec_tst;
