library verilog;
use verilog.vl_types.all;
entity counter4bit_vlg_vec_tst is
end counter4bit_vlg_vec_tst;
