library verilog;
use verilog.vl_types.all;
entity Divi_vlg_vec_tst is
end Divi_vlg_vec_tst;
