module lnx();
endmodule
