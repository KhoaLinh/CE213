library verilog;
use verilog.vl_types.all;
entity ControllerDecoder_vlg_vec_tst is
end ControllerDecoder_vlg_vec_tst;
