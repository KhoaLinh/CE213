library verilog;
use verilog.vl_types.all;
entity Lab2_CE221_vlg_vec_tst is
end Lab2_CE221_vlg_vec_tst;
