library verilog;
use verilog.vl_types.all;
entity SquareRoot_vlg_vec_tst is
end SquareRoot_vlg_vec_tst;
