library verilog;
use verilog.vl_types.all;
entity CAS8bit_vlg_vec_tst is
end CAS8bit_vlg_vec_tst;
