library verilog;
use verilog.vl_types.all;
entity counter8bit_parameter_vlg_vec_tst is
end counter8bit_parameter_vlg_vec_tst;
