library verilog;
use verilog.vl_types.all;
entity Squareroot_vlg_vec_tst is
end Squareroot_vlg_vec_tst;
