library verilog;
use verilog.vl_types.all;
entity tb_selfchecking is
end tb_selfchecking;
