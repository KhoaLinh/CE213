library verilog;
use verilog.vl_types.all;
entity getSignal_vlg_vec_tst is
end getSignal_vlg_vec_tst;
