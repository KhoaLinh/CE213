library verilog;
use verilog.vl_types.all;
entity counter_4bit_vlg_vec_tst is
end counter_4bit_vlg_vec_tst;
