library verilog;
use verilog.vl_types.all;
entity test_Squareroot_vlg_vec_tst is
end test_Squareroot_vlg_vec_tst;
