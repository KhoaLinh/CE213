library verilog;
use verilog.vl_types.all;
entity NextStageLogic_vlg_vec_tst is
end NextStageLogic_vlg_vec_tst;
