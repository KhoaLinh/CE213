library verilog;
use verilog.vl_types.all;
entity CAS17bit_vlg_vec_tst is
end CAS17bit_vlg_vec_tst;
