library verilog;
use verilog.vl_types.all;
entity lpm_counter_8bit_vlg_vec_tst is
end lpm_counter_8bit_vlg_vec_tst;
