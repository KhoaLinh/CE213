library verilog;
use verilog.vl_types.all;
entity C1_vlg_vec_tst is
end C1_vlg_vec_tst;
