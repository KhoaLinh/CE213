library verilog;
use verilog.vl_types.all;
entity testCounter is
end testCounter;
