library verilog;
use verilog.vl_types.all;
entity Controller_Decoder_vlg_vec_tst is
end Controller_Decoder_vlg_vec_tst;
