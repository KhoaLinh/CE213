library verilog;
use verilog.vl_types.all;
entity d_ff_struct_vlg_check_tst is
    port(
        q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end d_ff_struct_vlg_check_tst;
