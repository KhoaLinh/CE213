module MUXTRI6D(IN0, IN1, IN2, IN3, IN4, IN5, OUT, SEL);
input [15:0]IN0, IN1, IN2, IN3, IN4, IN5;
output [15:0]OUT;
input  SEL;

wire [15:0] OUT0, OUT1, OUT2, OUT3, OUT4, OUT;

MUXTRI MUXTRI0(IN0, IN1, SEL, OUT0);
MUXTRI MUXTRI1(IN2, IN3, SEL, OUT1);
MUXTRI MUXTRI2(IN4, IN5, SEL, OUT2);
MUXTRI MUXTRI3(OUT0, OUT1, SEL, OUT3);
MUXTRI MUXTRI4(OUT2, OUT3, SEL, OUT4);
MUXTRI MUXTRI5(OUT3, OUT4, SEL, OUT);



endmodule
