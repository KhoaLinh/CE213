library verilog;
use verilog.vl_types.all;
entity tb_lnx is
end tb_lnx;
