library verilog;
use verilog.vl_types.all;
entity clock_1s_vlg_vec_tst is
end clock_1s_vlg_vec_tst;
