library verilog;
use verilog.vl_types.all;
entity Multi_vlg_vec_tst is
end Multi_vlg_vec_tst;
