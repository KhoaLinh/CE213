library verilog;
use verilog.vl_types.all;
entity REG_vlg_vec_tst is
end REG_vlg_vec_tst;
