library verilog;
use verilog.vl_types.all;
entity test_Squareroot is
end test_Squareroot;
