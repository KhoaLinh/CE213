library verilog;
use verilog.vl_types.all;
entity Lab1_CE221_vlg_vec_tst is
end Lab1_CE221_vlg_vec_tst;
