library verilog;
use verilog.vl_types.all;
entity CounterCheck_vlg_check_tst is
    port(
        \OUT\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CounterCheck_vlg_check_tst;
