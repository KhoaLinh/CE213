library verilog;
use verilog.vl_types.all;
entity Counter12bit_vlg_vec_tst is
end Counter12bit_vlg_vec_tst;
