library verilog;
use verilog.vl_types.all;
entity counter_4bit_non_blocking_parameter_vlg_vec_tst is
end counter_4bit_non_blocking_parameter_vlg_vec_tst;
