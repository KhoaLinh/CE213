library verilog;
use verilog.vl_types.all;
entity C1_vlg_check_tst is
    port(
        Z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end C1_vlg_check_tst;
