library verilog;
use verilog.vl_types.all;
entity ROM_lab5_vlg_vec_tst is
end ROM_lab5_vlg_vec_tst;
