library verilog;
use verilog.vl_types.all;
entity CAS_vlg_vec_tst is
end CAS_vlg_vec_tst;
