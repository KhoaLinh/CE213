library verilog;
use verilog.vl_types.all;
entity twoDigitBCD_vlg_vec_tst is
end twoDigitBCD_vlg_vec_tst;
