library verilog;
use verilog.vl_types.all;
entity xorgate_vlg_vec_tst is
end xorgate_vlg_vec_tst;
